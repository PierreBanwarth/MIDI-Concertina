.title KiCad schematic
X1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 Net-_K15-Pad1_ NC_14 NC_15 NC_16 NC_17 NC_18 Net-_K?1-Pad1_ Net-_K14-Pad1_ NC_19 Net-_K1-Pad1_ Net-_K13-Pad1_ Net-_K2-Pad1_ Net-_K12-Pad1_ Net-_K3-Pad1_ Net-_K11-Pad1_ Net-_K4-Pad1_ Net-_K10-Pad1_ Net-_K5-Pad1_ Net-_K9-Pad1_ Net-_K6-Pad1_ Net-_K8-Pad1_ Net-_K7-Pad1_ Arduino_Pro_Mini
K?1 Net-_K?1-Pad1_ GND KEYSW
K1 Net-_K1-Pad1_ GND KEYSW
K2 Net-_K2-Pad1_ GND KEYSW
K3 Net-_K3-Pad1_ GND KEYSW
K4 Net-_K4-Pad1_ GND KEYSW
K5 Net-_K5-Pad1_ GND KEYSW
K6 Net-_K6-Pad1_ GND KEYSW
K7 Net-_K7-Pad1_ GND KEYSW
K8 Net-_K8-Pad1_ GND KEYSW
K9 Net-_K9-Pad1_ GND KEYSW
K10 Net-_K10-Pad1_ GND KEYSW
K11 Net-_K11-Pad1_ GND KEYSW
K12 Net-_K12-Pad1_ GND KEYSW
K13 Net-_K13-Pad1_ GND KEYSW
K14 Net-_K14-Pad1_ GND KEYSW
K15 Net-_K15-Pad1_ GND KEYSW
.end
